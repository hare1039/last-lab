module main ();
    
endmodule // main
